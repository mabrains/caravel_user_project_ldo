**.subckt ldo_v2
XM8 net2 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM9 net2 bg_out net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM10 net1 pos net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM11 net1 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM13 net3 vb GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM14 out net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12 
XM18 out vb GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12 
XM20 vb vb GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM24 ldo_out net5 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=800 m=800 
XM26 vb mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XC3 net1 net4 sky130_fd_pr__cap_mim_m3_1 W=60 L=60 MF=1 m=1
XR7 out net4 GND sky130_fd_pr__res_xhigh_po_0p69 L=4.5 mult=1 m=1
Vs VDD GND 2.3
Vt net6 GND 0
C2 net5 net6 5G m=1
L1 out net5 5G m=1
XR8 net7 ldo_out GND sky130_fd_pr__res_xhigh_po_0p69 L=24 mult=8 m=8
XR9 pos net7 GND sky130_fd_pr__res_xhigh_po_0p69 L=24 mult=3 m=3
XR12 net8 pos GND sky130_fd_pr__res_xhigh_po_0p69 L=24 mult=2 m=2
XR13 GND net8 GND sky130_fd_pr__res_xhigh_po_0p69 L=24 mult=4 m=4
XM1 inn mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM2 inp mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM3 bg_out mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XQ1 GND GND net10 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ5 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ6 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ7 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ9 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ11 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ13 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ15 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ17 GND GND net9 sky130_fd_pr__pnp_05v5_W0p68L0p68
XM7 net12 net12 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM12 net12 inp net11 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM21 mir inn net11 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM23 mir net12 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM15 net11 net13 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM25 net13 mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM16 net13 net13 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XC1 mir GND sky130_fd_pr__cap_mim_m3_1 W=16 L=16 MF=1 m=1
XR1 net14 inp GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=3 m=3
XR2 net10 inn GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=3 m=3
XR3 net16 net10 GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=1 m=1
XR10 net9 net14 GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=6 m=6
XR4 GND net15 GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=15 m=15
XR11 GND net16 GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=15 m=15
XR6 net15 net14 GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=1 m=1
XR5 net17 bg_out GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=1 m=1
XR14 GND net17 GND sky130_fd_pr__res_xhigh_po_0p69 L=27 mult=53 m=53
XM19 mir en VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
Ven en GND 2.3
XM4 net18 bg_out VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM5 net18 bg_out GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM6 VDD net18 inn GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
**** begin user architecture code


.param R=18k
R10 ldo_out GND {R}
IL ldo_out 0 PWL(0 0.1m 10u 0.1m 20u 10m 30u 10m)
*CL ldo_out gnd 10p
.lib /home/mustafa/mabrains/pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib_mod.spice tt




.nodeset v(inn)=1.2
.nodeset v(inp)=1.2
.nodeset v(mir)=1
.nodeset v(net13)=1
.nodeset v(bg_out)=1.1
.nodeset v(ldo_out)=1.8
.nodeset v(pos)=1.1
*.nodeset v(net3)=0.8
*.nodeset v(net1)=0.7
.nodeset v(net14)=0.9
*.nodeset v(net7)=0.75
.nodeset v(vb)=0.9

.option temp=27
*User_defined_functions
.control
define max(vector_name) (vecmax(vector_name))
define min(vector_name) (vecmin(vector_name))
.endc


*Temp_sweep
.control
alter IL 0
dc temp 85 0 -1
let temp_coeff=1000000*(max(ldo_out)-min(ldo_out))/85
print temp_coeff
plot v(ldo_out)
set wr_singlescale
set wr_vecnames
set appendwrite
.endc


.control
alter IL 0
*alter R10 1G
op
let iq =i(Vs)
print iq
*print all
set wr_singlescale
set wr_vecnames
set appendwrite
if v(ldo_out)>1
wrdata op_point_test v(ldo_out)
end
.endc



*Stability_Analysis
.control
alter IL 0
alter Vs AC =0
alter Vt AC=1
ac dec 10 1 1G
plot vdb(out)
plot (180/pi)*vp(out)
let ph= (180/pi)*vp(out)
meas ac pm FIND ph WHEN vdb(out)=0
.endc


*PSRR_Analysis
.control
alter IL 0
alter Vs AC =1
alter Vt AC=0
alter L1 0
alter C2 0
ac dec 10 1 1G
meas AC PSRR100 FIND vdb(ldo_out) AT=100
meas AC PSRR100k FIND vdb(ldo_out) AT=100k
plot vdb(ldo_out)
.endc




*supply_sweep
.control
alter IL 0
dc Vs 2.8 0 -0.01
plot vdd ldo_out
meas DC Vldo_Sup_2 FIND ldo_out AT=2
meas DC Vldo_nom FIND ldo_out AT=2.3
meas DC Vldo_Sup_2_8 FIND ldo_out AT=2.8
let line_reg = abs((Vldo_Sup_2_8-Vldo_Sup_2)/0.8)
print line_reg
meas DC vin WHEN v(ldo_out)=1.764
let dropout=vin-1.764
print dropout
set wr_singlescale
set wr_vecnames
set appendwrite
.endc





*Load_Reg_switches
*V1 c1 0 DC 0 PWL(0 5 20u 5 35u 0 50u 0 100u 0)
*V2 c2 0 DC 0 PWL(0 0 20u 0 35u 0 50u 5 100u 5)
*s1 ldo_out 2 c1 0 switch1 ON
*s2 ldo_out 3 c2 0 switch1 OFF
*.model switch1 sw vt=0.1 ron =0.1 roff =1G
*R1 2 0 18k
*R2 3 0 180

*.control
*alter R10 1G
*tran 0.1u 90u
*plot v(ldo_out) v(c1) v(c2)
*meas TRAN V_ldo_100u FIND v(ldo_out) AT=10u
*meas TRAN V_ldo_10m FIND v(ldo_out) AT=50u
*let load_reg= V_ldo_100u-V_ldo_10m
*print load_reg
*.endc


**Load_Transient
.control
alter IL 50u
alter R10 3600k
tran 0.1u 100u
meas TRAN V_ldo_100u FIND v(ldo_out) AT=5u
meas TRAN V_ldo_10m FIND v(ldo_out) AT=100u
let load_reg= V_ldo_100u-V_ldo_10m
let load_current =(-1*i(Vs)-131.8e-6)
print load_reg
plot load_current v(ldo_out)-1.8
.endc


**Transient
.control
alter R10 36k
alter @IL[PWL] = [ 0 0 10u 0 20u 0 30u 0 ]
alter @Vs[pulse] = [ 1 3 10u 10u 1u 100u 200u ]
alter IL 0
tran 0.1u 100u
plot vdd ldo_out
.endc

.control
alter R10 36k
alter @IL[PWL] = [ 0 0 10u 0 20u 0 30u 0 ]
alter @Vs[pulse] = [ 0 2.3 10u 0.1u 1u 100u 200u ]
tran 0.1u 100u
plot vdd ldo_out
.endc

.control
alter R10 36k
alter @IL[PWL] = [ 0 0 10u 0 20u 0 30u 0 ]
alter @Ven[pulse] = [ 0 2.3 10u 0.1u 1u 100u 200u ]
tran 0.1u 100u
*meas TRAN st_up_time when v(ldo_out)>1.782
plot en ldo_out
.endc





**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
** flattened .save nodes
.end
