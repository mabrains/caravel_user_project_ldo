**.subckt Error_Amp
**.ends
** flattened .save nodes
.end
